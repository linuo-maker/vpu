module xpu_vpu_pc_tn_vlsu_nan_checker(
    lane_data_has_nan，
    vlsu_lane_data，
    vlsu_lane_mew,
    vlsu_lane_strb
);
   // &Ports; @19
input   [127:0]  vlsu_lane_data;        
input   [1  :0]  vlsu_lane_mew;         
input   [15 :0]  vlsu_lane_strb;        
output           lane_data_has_nan;     

// &Regs; @20

// &Wires; @21
wire             bf16_has_nan;          
wire    [15 :0]  byte_ofp8_is_nan;      
wire    [1  :0]  dwrd_fp64_is_nan;      
wire             fp16_has_nan;          
wire             fp32_has_nan;          
wire             fp64_has_nan;          
wire    [7  :0]  half_bf16_is_nan;      
wire    [7  :0]  half_fp16_is_nan;      
wire    [127:0]  lane_data;             
wire             lane_data_has_nan;     
wire    [1  :0]  lane_mew;              
wire    [7  :0]  lane_split_data_byte0; 
wire    [7  :0]  lane_split_data_byte1; 
wire    [7  :0]  lane_split_data_byte10; 
wire    [7  :0]  lane_split_data_byte11; 
wire    [7  :0]  lane_split_data_byte12; 
wire    [7  :0]  lane_split_data_byte13; 
wire    [7  :0]  lane_split_data_byte14; 
wire    [7  :0]  lane_split_data_byte15; 
wire    [7  :0]  lane_split_data_byte2; 
wire    [7  :0]  lane_split_data_byte3; 
wire    [7  :0]  lane_split_data_byte4; 
wire    [7  :0]  lane_split_data_byte5; 
wire    [7  :0]  lane_split_data_byte6; 
wire    [7  :0]  lane_split_data_byte7; 
wire    [7  :0]  lane_split_data_byte8; 
wire    [7  :0]  lane_split_data_byte9; 
wire    [63 :0]  lane_split_data_dwrd0; 
wire    [63 :0]  lane_split_data_dwrd1; 
wire    [15 :0]  lane_split_data_half0; 
 wire    [15 :0]  lane_split_data_half1; 
wire    [15 :0]  lane_split_data_half2; 
wire    [15 :0]  lane_split_data_half3; 
wire    [15 :0]  lane_split_data_half4; 
wire    [15 :0]  lane_split_data_half5; 
wire    [15 :0]  lane_split_data_half6; 
wire    [15 :0]  lane_split_data_half7; 
wire    [31 :0]  lane_split_data_word0; 
wire    [31 :0]  lane_split_data_word1; 
wire    [31 :0]  lane_split_data_word2; 
wire    [31 :0]  lane_split_data_word3; 
wire    [15 :0]  lane_split_vld_byte;   
wire    [1  :0]  lane_split_vld_dwrd;   
wire    [7  :0]  lane_split_vld_half;   
wire    [3  :0]  lane_split_vld_word;   
wire    [15 :0]  lane_strb;             
wire             mew_bit8_sel;          
wire             mew_dwrd_sel;          
wire             mew_half_sel;          
wire             mew_word_sel;          
wire             ofp8_has_nan;          
wire    [127:0]  vlsu_lane_data;        
wire    [1  :0]  vlsu_lane_mew;         
wire    [15 :0]  vlsu_lane_strb;        
wire    [3  :0]  word_fp32_is_nan;      

//==========================================================================================||
//               I. Input                                                                   ||
//==========================================================================================||
assign lane_data[`XPU_VPU_PC_TN_LANE_VLEN-1:0]  = vlsu_lane_data[`XPU_VPU_PC_TN_LANE_VLEN-1:0];
assign lane_strb[`XPU_VPU_PC_TN_VLSU_ENUM-1:0]  = vlsu_lane_strb[`XPU_VPU_PC_TN_VLSU_ENUM-1:0];
assign lane_mew[1:0]                 = vlsu_lane_mew[1:0]               ;
//==========================================================================================||
//               II. Logic                                                                  ||
//==========================================================================================||
// -------------------------------------------------------------------------------------------
// II-1 Data split
// II-1.1 8-bit split
// &LoopGenBeg("zz",0,`XPU_VPU_PC_TN_LANE_VLEN/8-1); @35
// assign lane_split_data_bytezz[7:0]  = lane_data[zz*8+:8]; @36
// assign lane_split_vld_byte[zz]      = lane_strb[zz]; @37
assign lane_split_data_byte0[7:0]  = lane_data[0+:8];
assign lane_split_vld_byte[0]      = lane_strb[0];
assign lane_split_data_byte1[7:0]  = lane_data[8+:8];
assign lane_split_vld_byte[1]      = lane_strb[1];
assign lane_split_data_byte2[7:0]  = lane_data[16+:8];
assign lane_split_vld_byte[2]      = lane_strb[2];
assign lane_split_data_byte3[7:0]  = lane_data[24+:8];
assign lane_split_vld_byte[3]      = lane_strb[3];
assign lane_split_data_byte4[7:0]  = lane_data[32+:8];
assign lane_split_vld_byte[4]      = lane_strb[4];
assign lane_split_data_byte5[7:0]  = lane_data[40+:8];
assign lane_split_vld_byte[5]      = lane_strb[5];
assign lane_split_data_byte6[7:0]  = lane_data[48+:8];
assign lane_split_vld_byte[6]      = lane_strb[6];
assign lane_split_data_byte7[7:0]  = lane_data[56+:8];
assign lane_split_vld_byte[7]      = lane_strb[7];
assign lane_split_data_byte8[7:0]  = lane_data[64+:8];
assign lane_split_vld_byte[8]      = lane_strb[8];
assign lane_split_data_byte9[7:0]  = lane_data[72+:8];
assign lane_split_vld_byte[9]      = lane_strb[9];
assign lane_split_data_byte10[7:0]  = lane_data[80+:8];
assign lane_split_vld_byte[10]      = lane_strb[10];
assign lane_split_data_byte11[7:0]  = lane_data[88+:8];
assign lane_split_vld_byte[11]      = lane_strb[11];
assign lane_split_data_byte12[7:0]  = lane_data[96+:8];
assign lane_split_vld_byte[12]      = lane_strb[12];
assign lane_split_data_byte13[7:0]  = lane_data[104+:8];
assign lane_split_vld_byte[13]      = lane_strb[13];
assign lane_split_data_byte14[7:0]  = lane_data[112+:8];
assign lane_split_vld_byte[14]      = lane_strb[14];
assign lane_split_data_byte15[7:0]  = lane_data[120+:8];
assign lane_split_vld_byte[15]      = lane_strb[15];
// &LoopGenEnd; @38
// II-1.2 16-bit split
// &LoopGenBeg("zz",0,`XPU_VPU_PC_TN_LANE_VLEN/16-1); @40
// assign lane_split_data_halfzz[15:0] = lane_data[zz*16+:16]; @41
// assign lane_split_vld_half[zz]      = lane_strb[zz*2]; @42
assign lane_split_data_half0[15:0] = lane_data[0+:16];
assign lane_split_vld_half[0]      = lane_strb[0];
assign lane_split_data_half1[15:0] = lane_data[16+:16];
assign lane_split_vld_half[1]      = lane_strb[2];
assign lane_split_data_half2[15:0] = lane_data[32+:16];
assign lane_split_vld_half[2]      = lane_strb[4];
assign lane_split_data_half3[15:0] = lane_data[48+:16];
assign lane_split_vld_half[3]      = lane_strb[6];
assign lane_split_data_half4[15:0] = lane_data[64+:16];
assign lane_split_vld_half[4]      = lane_strb[8];
assign lane_split_data_half5[15:0] = lane_data[80+:16];
assign lane_split_vld_half[5]      = lane_strb[10];
assign lane_split_data_half6[15:0] = lane_data[96+:16];
assign lane_split_vld_half[6]      = lane_strb[12];
assign lane_split_data_half7[15:0] = lane_data[112+:16];
assign lane_split_vld_half[7]      = lane_strb[14];
// &LoopGenEnd; @43
// II-1.3 32-bit split
// &LoopGenBeg("zz",0,`XPU_VPU_PC_TN_LANE_VLEN/32-1); @45
// assign lane_split_data_wordzz[31:0] = lane_data[zz*32+:32]; @46
// assign lane_split_vld_word[zz]      = lane_strb[zz*4]; @47
assign lane_split_data_word0[31:0] = lane_data[0+:32];
assign lane_split_vld_word[0]      = lane_strb[0];
assign lane_split_data_word1[31:0] = lane_data[32+:32];
assign lane_split_vld_word[1]      = lane_strb[4];
assign lane_split_data_word2[31:0] = lane_data[64+:32];
assign lane_split_vld_word[2]      = lane_strb[8];
assign lane_split_data_word3[31:0] = lane_data[96+:32];
assign lane_split_vld_word[3]      = lane_strb[12];
// &LoopGenEnd; @48
// II-1.4 64-bit split
// &LoopGenBeg("zz",0,`XPU_VPU_PC_TN_LANE_VLEN/64-1); @50
// assign lane_split_data_dwrdzz[63:0] = lane_data[zz*64+:64]; @51
// assign lane_split_vld_dwrd[zz]      = lane_strb[zz*8]; @52
assign lane_split_data_dwrd0[63:0] = lane_data[0+:64];
assign lane_split_vld_dwrd[0]      = lane_strb[0];
assign lane_split_data_dwrd1[63:0] = lane_data[64+:64];
assign lane_split_vld_dwrd[1]      = lane_strb[8];
// &LoopGenEnd; @53
// II-1.5 mew select
assign mew_bit8_sel = ~(|lane_mew[1:0]);
assign mew_half_sel = ~lane_mew[1] &  lane_mew[0];
assign mew_word_sel =  lane_mew[1] & ~lane_mew[0];
assign mew_dwrd_sel = &lane_mew[1:0];
// -------------------------------------------------------------------------------------------
// II-2 Instance
// II-2.1 OFP8 NaN
// &LoopGenBeg("zz",0,`XPU_VPU_PC_TN_LANE_VLEN/8-1); @62
// &Instance("tn_vlsu_ofp8_nan_type","x_tn_vlsu_ofp8_nan_type_zz"); @63
// &Connect(.float_data(lane_split_data_bytezz[7:0])); @64
// &Connect(.is_nan(byte_ofp8_is_nan[zz])); @65
xpu_vpu_pc_tn_vlsu_ofp8_nan_type  x_tn_vlsu_ofp8_nan_type_0 (
  .float_data                 (lane_split_data_byte0[7:0]),
  .is_nan                     (byte_ofp8_is_nan[0]       )
);

xpu_vpu_pc_tn_vlsu_ofp8_nan_type  x_tn_vlsu_ofp8_nan_type_1 (
  .float_data                 (lane_split_data_byte1[7:0]),
  .is_nan                     (byte_ofp8_is_nan[1]       )
);

xpu_vpu_pc_tn_vlsu_ofp8_nan_type  x_tn_vlsu_ofp8_nan_type_2 (
  .float_data                 (lane_split_data_byte2[7:0]),
  .is_nan                     (byte_ofp8_is_nan[2]       )
);

xpu_vpu_pc_tn_vlsu_ofp8_nan_type  x_tn_vlsu_ofp8_nan_type_3 (
  .float_data                 (lane_split_data_byte3[7:0]),
  .is_nan                     (byte_ofp8_is_nan[3]       )
);

xpu_vpu_pc_tn_vlsu_ofp8_nan_type  x_tn_vlsu_ofp8_nan_type_4 (
  .float_data                 (lane_split_data_byte4[7:0]),
  .is_nan                     (byte_ofp8_is_nan[4]       )
);

xpu_vpu_pc_tn_vlsu_ofp8_nan_type  x_tn_vlsu_ofp8_nan_type_5 (
  .float_data                 (lane_split_data_byte5[7:0]),
  .is_nan                     (byte_ofp8_is_nan[5]       )
);

xpu_vpu_pc_tn_vlsu_ofp8_nan_type  x_tn_vlsu_ofp8_nan_type_6 (
  .float_data                 (lane_split_data_byte6[7:0]),
  .is_nan                     (byte_ofp8_is_nan[6]       )
);
xpu_vpu_pc_tn_vlsu_ofp8_nan_type  x_tn_vlsu_ofp8_nan_type_7 (
  .float_data                 (lane_split_data_byte7[7:0]),
  .is_nan                     (byte_ofp8_is_nan[7]       )
);

xpu_vpu_pc_tn_vlsu_ofp8_nan_type  x_tn_vlsu_ofp8_nan_type_8 (
  .float_data                 (lane_split_data_byte8[7:0]),
  .is_nan                     (byte_ofp8_is_nan[8]       )
);

xpu_vpu_pc_tn_vlsu_ofp8_nan_type  x_tn_vlsu_ofp8_nan_type_9 (
  .float_data                 (lane_split_data_byte9[7:0]),
  .is_nan                     (byte_ofp8_is_nan[9]       )
);

xpu_vpu_pc_tn_vlsu_ofp8_nan_type  x_tn_vlsu_ofp8_nan_type_10 (
  .float_data                  (lane_split_data_byte10[7:0]),
  .is_nan                      (byte_ofp8_is_nan[10]       )
);

xpu_vpu_pc_tn_vlsu_ofp8_nan_type  x_tn_vlsu_ofp8_nan_type_11 (
  .float_data                  (lane_split_data_byte11[7:0]),
  .is_nan                      (byte_ofp8_is_nan[11]       )
);

xpu_vpu_pc_tn_vlsu_ofp8_nan_type  x_tn_vlsu_ofp8_nan_type_12 (
  .float_data                  (lane_split_data_byte12[7:0]),
  .is_nan                      (byte_ofp8_is_nan[12]       )
);

xpu_vpu_pc_tn_vlsu_ofp8_nan_type  x_tn_vlsu_ofp8_nan_type_13 (
  .float_data                  (lane_split_data_byte13[7:0]),
  .is_nan                      (byte_ofp8_is_nan[13]       )
);

xpu_vpu_pc_tn_vlsu_ofp8_nan_type  x_tn_vlsu_ofp8_nan_type_14 (
  .float_data                  (lane_split_data_byte14[7:0]),
  .is_nan                      (byte_ofp8_is_nan[14]       )
);

xpu_vpu_pc_tn_vlsu_ofp8_nan_type  x_tn_vlsu_ofp8_nan_type_15 (
  .float_data                  (lane_split_data_byte15[7:0]),
  .is_nan                      (byte_ofp8_is_nan[15]       )
);

// &LoopGenEnd; @66
// II-2.2 BF16 NaN
// &LoopGenBeg("zz",0,`XPU_VPU_PC_TN_LANE_VLEN/16-1); @68
// &Instance("tn_vlsu_bf16_nan_type","x_tn_vlsu_bf16_nan_type_zz"); @69
// &Connect(.float_data(lane_split_data_halfzz[15:0])); @70
// &Connect(.is_nan(half_bf16_is_nan[zz])); @71
xpu_vpu_pc_tn_vlsu_bf16_nan_type  x_tn_vlsu_bf16_nan_type_0 (
  .float_data                  (lane_split_data_half0[15:0]),
  .is_nan                      (half_bf16_is_nan[0]        )
);

xpu_vpu_pc_tn_vlsu_bf16_nan_type  x_tn_vlsu_bf16_nan_type_1 (
  .float_data                  (lane_split_data_half1[15:0]),
  .is_nan                      (half_bf16_is_nan[1]        )
);

xpu_vpu_pc_tn_vlsu_bf16_nan_type  x_tn_vlsu_bf16_nan_type_2 (
  .float_data                  (lane_split_data_half2[15:0]),
  .is_nan                      (half_bf16_is_nan[2]        )
);

xpu_vpu_pc_tn_vlsu_bf16_nan_type  x_tn_vlsu_bf16_nan_type_3 (
  .float_data                  (lane_split_data_half3[15:0]),
  .is_nan                      (half_bf16_is_nan[3]        )
);

xpu_vpu_pc_tn_vlsu_bf16_nan_type  x_tn_vlsu_bf16_nan_type_4 (
  .float_data                  (lane_split_data_half4[15:0]),
  .is_nan                      (half_bf16_is_nan[4]        )
);

xpu_vpu_pc_tn_vlsu_bf16_nan_type  x_tn_vlsu_bf16_nan_type_5 (
  .float_data                  (lane_split_data_half5[15:0]),
  .is_nan                      (half_bf16_is_nan[5]        )
);

xpu_vpu_pc_tn_vlsu_bf16_nan_type  x_tn_vlsu_bf16_nan_type_6 (
  .float_data                  (lane_split_data_half6[15:0]),
  .is_nan                      (half_bf16_is_nan[6]        )
);

xpu_vpu_pc_tn_vlsu_bf16_nan_type  x_tn_vlsu_bf16_nan_type_7 (
  .float_data                  (lane_split_data_half7[15:0]),
  .is_nan                      (half_bf16_is_nan[7]        )
);

// &LoopGenEnd; @72
// II-2.3 IEEE754 FP16 NaN
// &LoopGenBeg("zz",0,`XPU_VPU_PC_TN_LANE_VLEN/16-1); @74
// &Instance('#(.EXPONENT_SIZE(5), .MANTISSA_SIZE(10))', "tn_vlsu_ieee754_nan_type", "x_tn_vl @75
// &Connect(.float_data(lane_split_data_halfzz[15:0])); @76
// &Connect(.is_nan(half_fp16_is_nan[zz])); @77
xpu_vpu_pc_tn_vlsu_ieee754_nan_type #(.EXPONENT_SIZE(5), .MANTISSA_SIZE(10)) x_tn_vlsu_ieee754_nan_type_fp16_0 (
  .float_data                  (lane_split_data_half0[15:0]),
  .is_nan                      (half_fp16_is_nan[0]        )
);

xpu_vpu_pc_tn_vlsu_ieee754_nan_type #(.EXPONENT_SIZE(5), .MANTISSA_SIZE(10)) x_tn_vlsu_ieee754_nan_type_fp16_1 (
  .float_data                  (lane_split_data_half1[15:0]),
  .is_nan                      (half_fp16_is_nan[1]        )
);

xpu_vpu_pc_tn_vlsu_ieee754_nan_type #(.EXPONENT_SIZE(5), .MANTISSA_SIZE(10)) x_tn_vlsu_ieee754_nan_type_fp16_2 (
  .float_data                  (lane_split_data_half2[15:0]),
  .is_nan                      (half_fp16_is_nan[2]        )
);

xpu_vpu_pc_tn_vlsu_ieee754_nan_type #(.EXPONENT_SIZE(5), .MANTISSA_SIZE(10)) x_tn_vlsu_ieee754_nan_type_fp16_3 (
  .float_data                  (lane_split_data_half3[15:0]),
  .is_nan                      (half_fp16_is_nan[3]        )
);

xpu_vpu_pc_tn_vlsu_ieee754_nan_type #(.EXPONENT_SIZE(5), .MANTISSA_SIZE(10)) x_tn_vlsu_ieee754_nan_type_fp16_4 (
  .float_data                  (lane_split_data_half4[15:0]),
  .is_nan                      (half_fp16_is_nan[4]        )
);

xpu_vpu_pc_tn_vlsu_ieee754_nan_type #(.EXPONENT_SIZE(5), .MANTISSA_SIZE(10)) x_tn_vlsu_ieee754_nan_type_fp16_5 (
  .float_data                  (lane_split_data_half5[15:0]),
  .is_nan                      (half_fp16_is_nan[5]        )
);

xpu_vpu_pc_tn_vlsu_ieee754_nan_type #(.EXPONENT_SIZE(5), .MANTISSA_SIZE(10)) x_tn_vlsu_ieee754_nan_type_fp16_6 (
  .float_data                  (lane_split_data_half6[15:0]),
  .is_nan                      (half_fp16_is_nan[6]        )
);

xpu_vpu_pc_tn_vlsu_ieee754_nan_type #(.EXPONENT_SIZE(5), .MANTISSA_SIZE(10)) x_tn_vlsu_ieee754_nan_type_fp16_7 (
  .float_data                  (lane_split_data_half7[15:0]),
  .is_nan                      (half_fp16_is_nan[7]        )
);

// &LoopGenEnd; @78
// II-2.4 IEEE754 FP32 NaN
// &LoopGenBeg("zz",0,`XPU_VPU_PC_TN_LANE_VLEN/32-1); @80
// &Instance('#(.EXPONENT_SIZE(8), .MANTISSA_SIZE(23))', "tn_vlsu_ieee754_nan_type", "x_tn_vl @81
// &Connect(.float_data(lane_split_data_wordzz[31:0])); @82
// &Connect(.is_nan(word_fp32_is_nan[zz])); @83
xpu_vpu_pc_tn_vlsu_ieee754_nan_type #(.EXPONENT_SIZE(8), .MANTISSA_SIZE(23)) x_tn_vlsu_ieee754_nan_type_fp32_0 (
  .float_data                  (lane_split_data_word0[31:0]),
  .is_nan                      (word_fp32_is_nan[0]        )
);

xpu_vpu_pc_tn_vlsu_ieee754_nan_type #(.EXPONENT_SIZE(8), .MANTISSA_SIZE(23)) x_tn_vlsu_ieee754_nan_type_fp32_1 (
  .float_data                  (lane_split_data_word1[31:0]),
  .is_nan                      (word_fp32_is_nan[1]        )
);

xpu_vpu_pc_tn_vlsu_ieee754_nan_type #(.EXPONENT_SIZE(8), .MANTISSA_SIZE(23)) x_tn_vlsu_ieee754_nan_type_fp32_2 (
  .float_data                  (lane_split_data_word2[31:0]),
  .is_nan                      (word_fp32_is_nan[2]        )
);

xpu_vpu_pc_tn_vlsu_ieee754_nan_type #(.EXPONENT_SIZE(8), .MANTISSA_SIZE(23)) x_tn_vlsu_ieee754_nan_type_fp32_3 (
  .float_data                  (lane_split_data_word3[31:0]),
  .is_nan                      (word_fp32_is_nan[3]        )
);

// &LoopGenEnd; @84
// II-2.5 IEEE754 FP64 NaN
// &LoopGenBeg("zz",0,`XPU_VPU_PC_TN_LANE_VLEN/64-1); @86
// &Instance('#(.EXPONENT_SIZE(11), .MANTISSA_SIZE(52))', "tn_vlsu_ieee754_nan_type", "x_tn_v @87
// &Connect(.float_data(lane_split_data_dwrdzz[63:0])); @88
// &Connect(.is_nan(dwrd_fp64_is_nan[zz])); @89
xpu_vpu_pc_tn_vlsu_ieee754_nan_type #(.EXPONENT_SIZE(11), .MANTISSA_SIZE(52)) x_tn_vlsu_ieee754_nan_type_fp64_0 (
  .float_data                  (lane_split_data_dwrd0[63:0]),
  .is_nan                      (dwrd_fp64_is_nan[0]        )
);

xpu_vpu_pc_tn_vlsu_ieee754_nan_type #(.EXPONENT_SIZE(11), .MANTISSA_SIZE(52)) x_tn_vlsu_ieee754_nan_type_fp64_1 (
  .float_data                  (lane_split_data_dwrd1[63:0]),
  .is_nan                      (dwrd_fp64_is_nan[1]        )
);

// &LoopGenEnd; @90
// -------------------------------------------------------------------------------------------
// II-3 Result comb
assign ofp8_has_nan = |(byte_ofp8_is_nan[`XPU_VPU_PC_TN_LANE_VLEN/8-1:0] 
                    & lane_split_vld_byte[`XPU_VPU_PC_TN_LANE_VLEN/8-1:0]);
assign bf16_has_nan = |(half_bf16_is_nan[`XPU_VPU_PC_TN_LANE_VLEN/16-1:0] 
                    & lane_split_vld_half[`XPU_VPU_PC_TN_LANE_VLEN/16-1:0]);
assign fp16_has_nan = |(half_fp16_is_nan[`XPU_VPU_PC_TN_LANE_VLEN/16-1:0] 
                    & lane_split_vld_half[`XPU_VPU_PC_TN_LANE_VLEN/16-1:0]);
assign fp32_has_nan = |(word_fp32_is_nan[`XPU_VPU_PC_TN_LANE_VLEN/32-1:0] 
                    & lane_split_vld_word[`XPU_VPU_PC_TN_LANE_VLEN/32-1:0]);
assign fp64_has_nan = |(dwrd_fp64_is_nan[`XPU_VPU_PC_TN_LANE_VLEN/64-1:0] 
                    & lane_split_vld_dwrd[`XPU_VPU_PC_TN_LANE_VLEN/64-1:0]);
//==========================================================================================||
//              III. Output                                                                 ||
//==========================================================================================||
assign lane_data_has_nan            = ofp8_has_nan & mew_bit8_sel
                                    | bf16_has_nan & mew_half_sel
                                    | fp16_has_nan & mew_half_sel
                                    | fp32_has_nan & mew_word_sel
                                    | fp64_has_nan & mew_dwrd_sel;

// &ModuleEnd; @112
endmodule
